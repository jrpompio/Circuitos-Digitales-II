module test (/*AUTOARG*/);

