module ejemplomode(/*AUTOARG*/
   // Outputs
   B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, B11, B12, B13, B14, B15,
   B16, B17, B18, B19, B20, B21, B22, B23, B24, B25, B26, B27, B28,
   B29, B30, B31, B32, B33, B34, B35, B36, B37, B38, B39, B40, B41,
   // Inputs
   A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15,
   A16, A17, A18, A19, A20, A21
   );
   /*AUTOINPUT*/
	 input wire A1;
	 input wire A2;
	 input wire A3;
	 input wire A4;
	 input wire A5;
	 input wire A6;
	 input wire A7;
	 input wire A8;
	 input wire A9;
	 input wire A10;
	 input wire A11;
	 input wire A12;
	 input wire A13;
	 input wire A14;
	 input wire A15;
	 input wire A16;
	 input wire A17;
	 input wire A18;
	 input wire A19;
	 input wire A20;
	 input wire A21;
   /*AUTOOUTPUT*/
   output reg B1;
   output reg B2;
   output reg B3;
   output reg B4;
   output reg B5;
   output reg B6;
   output reg B7;
   output reg B8;
   output reg B9;
   output reg B10;
   output reg B11;
   output reg B12;
   output reg B13;
   output reg B14;
   output reg B15;
   output reg B16;
   output reg B17;
   output reg B18;
   output reg B19;
   output reg B20;
   output reg B21;
   output reg B22;
   output reg B23;
   output reg B24;
   output reg B25;
   output reg B26;
   output reg B27;
   output reg B28;
   output reg B29;
   output reg B30;
   output reg B31;
   output reg B32;
   output reg B33;
   output reg B34;
   output reg B35;
   output reg B36;
   output reg B37;
   output reg B38;
   output reg B39;
   output reg B40;
   output reg B41;

ejemplomode instancia (/*AUTOINST*/
		       // Outputs
		       .B1		(B1),
		       .B2		(B2),
		       .B3		(B3),
		       .B4		(B4),
		       .B5		(B5),
		       .B6		(B6),
		       .B7		(B7),
		       .B8		(B8),
		       .B9		(B9),
		       .B10		(B10),
		       .B11		(B11),
		       .B12		(B12),
		       .B13		(B13),
		       .B14		(B14),
		       .B15		(B15),
		       .B16		(B16),
		       .B17		(B17),
		       .B18		(B18),
		       .B19		(B19),
		       .B20		(B20),
		       .B21		(B21),
		       .B22		(B22),
		       .B23		(B23),
		       .B24		(B24),
		       .B25		(B25),
		       .B26		(B26),
		       .B27		(B27),
		       .B28		(B28),
		       .B29		(B29),
		       .B30		(B30),
		       .B31		(B31),
		       .B32		(B32),
		       .B33		(B33),
		       .B34		(B34),
		       .B35		(B35),
		       .B36		(B36),
		       .B37		(B37),
		       .B38		(B38),
		       .B39		(B39),
		       .B40		(B40),
		       .B41		(B41),
		       // Inputs
		       .A1		(A1),
		       .A2		(A2),
		       .A3		(A3),
		       .A4		(A4),
		       .A5		(A5),
		       .A6		(A6),
		       .A7		(A7),
		       .A8		(A8),
		       .A9		(A9),
		       .A10		(A10),
		       .A11		(A11),
		       .A12		(A12),
		       .A13		(A13),
		       .A14		(A14),
		       .A15		(A15),
		       .A16		(A16),
		       .A17		(A17),
		       .A18		(A18),
		       .A19		(A19),
		       .A20		(A20),
		       .A21		(A21));

endmodule



